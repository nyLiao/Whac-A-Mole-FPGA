module wam_led (
    input wire [7:0] sw,
    output reg [3:0] ld
    );

    

endmodule // wam_led
